`include "configs.v"

module ID_Stage_Reg(
  input clk, rst,
  input[`ADDRESS_LEN - 1:0] pc_in,
  output reg[`ADDRESS_LEN - 1:0] pc
);
  
  
endmodule