`include "configs.v"

module Val2_Generator(
  input [31:0] Val_Rm,
  input [11:0] Shift_operand,
  input imm, is_mem,
  output [31:0] Val2
);

  

endmodule