`include "configs.v"

module Instruction_Memory(output reg[`WORD_LEN - 1 : 0] instruction, input[`ADDRESS_LEN - 1 : 0] address);
  reg [`WORD_LEN-1:0] regs[0:`MEMORY_SIZE-1];
  wire[`ADDRESS_LEN - 3 : 0] aligned_address = address[`WORD_LEN - 1:2];
  
  initial begin
    //regs[0] = 32'b00001000000000000000000001100100;// jmp 100
    regs[0] = 32'b00000000000000000000000000000000;// nop;
    regs[1] = 32'b1110_00_1_1101_0_0000_0000_000000010100; //MOVR0 ,#20 //R0 = 20
    regs[2] = 32'b1110_00_1_1101_0_0000_0001_101000000001; //MOVR1 ,#4096//R1 = 4096
    regs[3] = 32'b1110_00_1_1101_0_0000_0010_000100000011; //MOVR2 ,#0xC0000000//R2 = -1073741824
    regs[4] = 32'b1110_00_0_0100_1_0010_0011_000000000010; //ADDSR3 ,R2,R2//R3 = -2147483648 
    regs[5] = 32'b1110_00_0_0101_0_0000_0100_000000000000; //ADCR4 ,R0,R0//R4 = 41
    regs[6] = 32'b1110_00_0_0010_0_0100_0101_000100000100; //SUBR5 ,R4,R4,LSL #2//R5 = -123
    regs[7] = 32'b1110_00_0_0110_0_0000_0110_000010100000; //SBCR6 ,R0,R0,LSR #1//R6 = 10
    regs[8] = 32'b1110_00_0_1100_0_0101_0111_000101000010; //ORRR7 ,R5,R2,ASR #2//R7 = -123
    regs[9] = 32'b1110_00_0_0000_0_0111_1000_000000000011; //ANDR8 ,R7,R3//R8 = -2147483648
    regs[10] = 32'b1110_00_0_1111_0_0000_1001_000000000110; //MVNR9 ,R6//R9 = -11
    regs[11] = 32'b1110_00_0_0001_0_0100_1010_000000000101; //EORR10,R4,R5//R10 = -84
    regs[12] = 32'b1110_00_0_1010_1_1000_0000_000000000110; //CMPR8 ,R6
    regs[13] = 32'b0001_00_0_0100_0_0001_0001_000000000001; //ADDNER1 ,R1,R1//R1 = 8192
    regs[14] = 32'b1110_00_0_1000_1_1001_0000_000000001000; //TSTR9 ,R8
    regs[15] = 32'b0000_00_0_0100_0_0010_0010_000000000010; //ADDEQR2 ,R2,R2   //R2 = -1073741824
    regs[16] = 32'b1110_00_1_1101_0_0000_0000_101100000001; //MOVR0 ,#1024//R0 = 1024
    regs[17] = 32'b1110_01_0_0100_0_0000_0001_000000000000; //STRR1 ,[R0],#0//MEM[1024] = 8192
    regs[18] = 32'b1110_01_0_0100_1_0000_1011_000000000000; //LDRR11,[R0],#0//R11 = 8192
    regs[19] = 32'b1110_01_0_0100_0_0000_0010_000000000100; //STRR2 ,[R0],#4//MEM[1028] = -1073741824
    regs[20] = 32'b1110_01_0_0100_0_0000_0011_000000001000; //STRR3 ,[R0],#8//MEM[1032] = -2147483648
    regs[21] = 32'b1110_01_0_0100_0_0000_0100_000000001101; //STRR4 ,[R0],#13//MEM[1036] = 41
    regs[22] = 32'b1110_01_0_0100_0_0000_0101_000000010000; //STRR5 ,[R0],#16//MEM[1040] = -123
    regs[23] = 32'b1110_01_0_0100_0_0000_0110_000000010100; //STRR6,[R0],#20//MEM[1044] = 10
    regs[24] = 32'b1110_01_0_0100_1_0000_1010_000000000100; //LDRR10,[R0],#4//R10 = -1073741824
    regs[25] = 32'b1110_01_0_0100_0_0000_0111_000000011000; //STRR7 ,[R0],#24//MEM[1048] = -123
    regs[26] = 32'b1110_00_1_1101_0_0000_0001_000000000100; //MOVR1 ,#4//R1 = 4
    regs[27] = 32'b1110_00_1_1101_0_0000_0010_000000000000; //MOVR2 ,#0//R2 = 0
    regs[28] = 32'b1110_00_1_1101_0_0000_0011_000000000000; //MOVR3 ,#0//R3 = 0
    regs[29] = 32'b1110_00_0_0100_0_0000_0100_000100000011; //ADDR4 ,R0,R3,LSL #2
    regs[30] = 32'b1110_01_0_0100_1_0100_0101_000000000000; //LDRR5 ,[R4],#0
    regs[31] = 32'b1110_01_0_0100_1_0100_0110_000000000100; //LDRR6 ,[R4],#4
    regs[32] = 32'b1110_00_0_1010_1_0101_0000_000000000110; //CMPR5 ,R6
    regs[33] = 32'b1100_01_0_0100_0_0100_0110_000000000000; //STRGTR6 ,[R4],#0
    regs[34] = 32'b1100_01_0_0100_0_0100_0101_000000000100; //STRGTR5 ,[R4],#4
    regs[35] = 32'b1110_00_1_0100_0_0011_0011_000000000001; //ADDR3 ,R3,#1
    regs[36] = 32'b1110_00_1_1010_1_0011_0000_000000000011; //CMPR3 ,#3
    regs[37] = 32'b1011_10_1_0_111111111111111111110111  ; //BLT#-9
    regs[38] = 32'b1110_00_1_0100_0_0010_0010_000000000001; //ADDR2 ,R2,#1
    regs[39] = 32'b1110_00_0_1010_1_0010_0000_000000000001;//CMPR2 ,R1
    regs[40] = 32'b1011_10_1_0_111111111111111111110011  ;//BLT#-13
    regs[41] = 32'b1110_01_0_0100_1_0000_0001_000000000000;//LDRR1 ,[R0],#0//R1 = -2147483648
    regs[42] = 32'b1110_01_0_0100_1_0000_0010_000000000100;//LDRR2 ,[R0],#4//R2 = -1073741824
    regs[43] = 32'b1110_01_0_0100_1_0000_0011_000000001000;//STRR3 ,[R0],#8//R3 = 41
    regs[44] = 32'b1110_01_0_0100_1_0000_0100_000000001100;//STRR4 ,[R0],#12//R4 = 8192
    regs[45] = 32'b1110_01_0_0100_1_0000_0101_000000010000;//STRR5 ,[R0],#16//R5= -123
    regs[46] = 32'b1110_01_0_0100_1_0000_0110_000000010100;//STRR6 ,[R0],#20//R4 = 10
    regs[47] = 32'b1110_10_1_0_111111111111111111111111  ;//B#-1
    regs[48] = 32'b00000000000000000000000000000000;// nop;
    regs[49] = 32'b00000000000000000000000000000000;// nop;
    regs[50] = 32'b00000000000000000000000000000000;// nop;
    regs[51] = 32'b00000000000000000000000000000000;// nop;
    regs[52] = 32'b00000000000000000000000000000000;// nop;
    regs[53] = 32'b00000000000000000000000000000000;// nop;
    regs[54] = 32'b00000000000000000000000000000000;// nop;
    regs[55] = 32'b00000000000000000000000000000000;// nop;
    regs[56] = 32'b00000000000000000000000000000000;// nop;
  end

  always @(address) begin
    instruction = regs[aligned_address];
    //if(aligned_address < 40)
      //$display("CLK%d:--%b--", aligned_address, regs[aligned_address]);
  end

endmodule